LavaStatus=0
   XM    �          �  e 
    �  e  `   <   ( rW�F���     1< 2    V   G         [ 2V      ,2j   j   .2�   h   2         N i o s   I I   p r o c e s s o r   f o r   t h e   g a m e - 2 0 2 1 1 1 0 2 . z i p m s e d g e . e x e h t t p s : / / m o o d l e . e p f l . c h / m o d / f o l d e r / d o w n l o a d _ f o l d e r . p h p h t t p s : / / m o o d l e . e p f l . c h / m o d / f o l d e r / v i e w . p h p ? i d = 9 6 5 9 5 5 x$�